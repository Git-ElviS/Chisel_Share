module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  wire  _T = state_3 ^ state_2; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_2 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_3 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BasicRotate(
  input   clock,
  input   reset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  shiftAmount_prng_clock; // @[PRNG.scala 91:22]
  wire  shiftAmount_prng_reset; // @[PRNG.scala 91:22]
  wire  shiftAmount_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  shiftAmount_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  shiftAmount_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  shiftAmount_prng_io_out_3; // @[PRNG.scala 91:22]
  wire [3:0] shiftAmount = {shiftAmount_prng_io_out_3,shiftAmount_prng_io_out_2,shiftAmount_prng_io_out_1,
    shiftAmount_prng_io_out_0}; // @[PRNG.scala 95:17]
  reg [3:0] ctr; // @[UIntOps.scala 118:20]
  wire [2:0] _rotL_T_7 = shiftAmount[0] ? 3'h2 : 3'h1; // @[UIntOps.scala 120:33]
  wire [2:0] _rotL_T_10 = {_rotL_T_7[0],_rotL_T_7[2:1]}; // @[UIntOps.scala 120:33]
  wire [2:0] _rotL_T_11 = shiftAmount[1] ? _rotL_T_10 : _rotL_T_7; // @[UIntOps.scala 120:33]
  wire [2:0] _rotL_T_14 = {_rotL_T_11[1:0],_rotL_T_11[2]}; // @[UIntOps.scala 120:33]
  wire [2:0] _rotL_T_15 = shiftAmount[2] ? _rotL_T_14 : _rotL_T_11; // @[UIntOps.scala 120:33]
  wire [2:0] _rotL_T_18 = {_rotL_T_15[0],_rotL_T_15[2:1]}; // @[UIntOps.scala 120:33]
  wire [2:0] rotL = shiftAmount[3] ? _rotL_T_18 : _rotL_T_15; // @[UIntOps.scala 120:33]
  wire [2:0] _rotR_T_6 = shiftAmount[0] ? 3'h4 : 3'h1; // @[UIntOps.scala 121:34]
  wire [2:0] _rotR_T_9 = {_rotR_T_6[1:0],_rotR_T_6[2]}; // @[UIntOps.scala 121:34]
  wire [2:0] _rotR_T_10 = shiftAmount[1] ? _rotR_T_9 : _rotR_T_6; // @[UIntOps.scala 121:34]
  wire [2:0] _rotR_T_13 = {_rotR_T_10[0],_rotR_T_10[2:1]}; // @[UIntOps.scala 121:34]
  wire [2:0] _rotR_T_14 = shiftAmount[2] ? _rotR_T_13 : _rotR_T_10; // @[UIntOps.scala 121:34]
  wire [2:0] _rotR_T_17 = {_rotR_T_14[1:0],_rotR_T_14[2]}; // @[UIntOps.scala 121:34]
  wire [2:0] rotR = shiftAmount[3] ? _rotR_T_17 : _rotR_T_14; // @[UIntOps.scala 121:34]
  wire  _T_1 = ~reset; // @[UIntOps.scala 123:9]
  wire [3:0] _GEN_1 = shiftAmount % 4'h3; // @[UIntOps.scala 125:22]
  wire  _T_5 = 2'h0 == _GEN_1[1:0] | 2'h3 == _GEN_1[1:0]; // @[UIntOps.scala 125:29]
  wire  _T_14 = 2'h1 == _GEN_1[1:0]; // @[UIntOps.scala 125:29]
  wire  _T_23 = 2'h2 == _GEN_1[1:0]; // @[UIntOps.scala 125:29]
  wire [3:0] _ctr_T_1 = ctr + 4'h1; // @[UIntOps.scala 140:14]
  wire  _T_32 = ctr == 4'hf; // @[UIntOps.scala 142:12]
  wire  _GEN_0 = _T_5 & _T_1; // @[UIntOps.scala 127:13]
  wire  _GEN_6 = ~_T_5; // @[UIntOps.scala 131:13]
  wire  _GEN_8 = ~_T_5 & _T_14 & _T_1; // @[UIntOps.scala 131:13]
  wire  _GEN_24 = _GEN_6 & ~_T_14 & _T_23 & _T_1; // @[UIntOps.scala 135:13]
  MaxPeriodFibonacciLFSR shiftAmount_prng ( // @[PRNG.scala 91:22]
    .clock(shiftAmount_prng_clock),
    .reset(shiftAmount_prng_reset),
    .io_out_0(shiftAmount_prng_io_out_0),
    .io_out_1(shiftAmount_prng_io_out_1),
    .io_out_2(shiftAmount_prng_io_out_2),
    .io_out_3(shiftAmount_prng_io_out_3)
  );
  assign shiftAmount_prng_clock = clock;
  assign shiftAmount_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[UIntOps.scala 118:20]
      ctr <= 4'h0; // @[UIntOps.scala 118:20]
    end else begin
      ctr <= _ctr_T_1; // @[UIntOps.scala 140:7]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"Shift amount: %d rotateLeft:%b rotateRight:%b\n",shiftAmount,rotL,rotR); // @[UIntOps.scala 123:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_5 & _T_1 & ~(rotL == 3'h1)) begin
          $fatal; // @[UIntOps.scala 127:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_5 & _T_1 & ~(rotL == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UIntOps.scala:127 assert(rotL === \"b001\".U)\n"); // @[UIntOps.scala 127:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_0 & ~(rotR == 3'h1)) begin
          $fatal; // @[UIntOps.scala 128:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_0 & ~(rotR == 3'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UIntOps.scala:128 assert(rotR === \"b001\".U)\n"); // @[UIntOps.scala 128:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_5 & _T_14 & _T_1 & ~(rotL == 3'h2)) begin
          $fatal; // @[UIntOps.scala 131:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_5 & _T_14 & _T_1 & ~(rotL == 3'h2)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UIntOps.scala:131 assert(rotL === \"b010\".U)\n"); // @[UIntOps.scala 131:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_8 & ~(rotR == 3'h4)) begin
          $fatal; // @[UIntOps.scala 132:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_8 & ~(rotR == 3'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UIntOps.scala:132 assert(rotR === \"b100\".U)\n"); // @[UIntOps.scala 132:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_6 & ~_T_14 & _T_23 & _T_1 & ~(rotL == 3'h4)) begin
          $fatal; // @[UIntOps.scala 135:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_6 & ~_T_14 & _T_23 & _T_1 & ~(rotL == 3'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UIntOps.scala:135 assert(rotL === \"b100\".U)\n"); // @[UIntOps.scala 135:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_24 & ~(rotR == 3'h2)) begin
          $fatal; // @[UIntOps.scala 136:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_24 & ~(rotR == 3'h2)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UIntOps.scala:136 assert(rotR === \"b010\".U)\n"); // @[UIntOps.scala 136:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_32 & _T_1) begin
          $finish; // @[UIntOps.scala 143:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctr = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
