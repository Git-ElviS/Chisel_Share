module PassthroughModule(
  input  [31:0] io_in,
  output [31:0] io_out
);
  assign io_out = io_in; // @[Util.scala 19:10]
endmodule
module BidirectionalTester3DTabulate(
  input   clock,
  input   reset
);
  wire [31:0] PassthroughModule_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_1_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_1_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_2_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_2_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_3_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_3_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_4_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_4_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_5_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_5_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_6_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_6_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_7_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_7_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_8_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_8_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_9_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_9_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_10_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_10_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_11_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_11_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_12_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_12_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_13_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_13_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_14_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_14_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_15_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_15_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_16_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_16_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_17_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_17_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_18_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_18_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_19_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_19_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_20_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_20_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_21_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_21_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_22_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_22_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_23_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_23_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_24_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_24_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_25_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_25_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_26_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_26_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_27_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_27_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_28_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_28_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_29_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_29_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_30_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_30_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_31_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_31_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_32_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_32_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_33_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_33_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_34_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_34_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_35_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_35_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_36_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_36_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_37_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_37_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_38_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_38_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_39_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_39_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_40_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_40_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_41_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_41_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_42_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_42_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_43_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_43_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_44_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_44_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_45_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_45_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_46_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_46_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_47_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_47_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_48_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_48_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_49_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_49_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_50_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_50_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_51_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_51_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_52_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_52_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_53_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_53_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_54_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_54_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_55_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_55_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_56_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_56_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_57_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_57_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_58_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_58_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_59_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_59_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_60_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_60_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_61_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_61_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_62_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_62_io_out; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_63_io_in; // @[Vec.scala 225:30]
  wire [31:0] PassthroughModule_63_io_out; // @[Vec.scala 225:30]
  wire  _T_2 = ~reset; // @[Vec.scala 227:13]
  PassthroughModule PassthroughModule ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_io_in),
    .io_out(PassthroughModule_io_out)
  );
  PassthroughModule PassthroughModule_1 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_1_io_in),
    .io_out(PassthroughModule_1_io_out)
  );
  PassthroughModule PassthroughModule_2 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_2_io_in),
    .io_out(PassthroughModule_2_io_out)
  );
  PassthroughModule PassthroughModule_3 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_3_io_in),
    .io_out(PassthroughModule_3_io_out)
  );
  PassthroughModule PassthroughModule_4 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_4_io_in),
    .io_out(PassthroughModule_4_io_out)
  );
  PassthroughModule PassthroughModule_5 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_5_io_in),
    .io_out(PassthroughModule_5_io_out)
  );
  PassthroughModule PassthroughModule_6 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_6_io_in),
    .io_out(PassthroughModule_6_io_out)
  );
  PassthroughModule PassthroughModule_7 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_7_io_in),
    .io_out(PassthroughModule_7_io_out)
  );
  PassthroughModule PassthroughModule_8 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_8_io_in),
    .io_out(PassthroughModule_8_io_out)
  );
  PassthroughModule PassthroughModule_9 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_9_io_in),
    .io_out(PassthroughModule_9_io_out)
  );
  PassthroughModule PassthroughModule_10 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_10_io_in),
    .io_out(PassthroughModule_10_io_out)
  );
  PassthroughModule PassthroughModule_11 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_11_io_in),
    .io_out(PassthroughModule_11_io_out)
  );
  PassthroughModule PassthroughModule_12 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_12_io_in),
    .io_out(PassthroughModule_12_io_out)
  );
  PassthroughModule PassthroughModule_13 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_13_io_in),
    .io_out(PassthroughModule_13_io_out)
  );
  PassthroughModule PassthroughModule_14 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_14_io_in),
    .io_out(PassthroughModule_14_io_out)
  );
  PassthroughModule PassthroughModule_15 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_15_io_in),
    .io_out(PassthroughModule_15_io_out)
  );
  PassthroughModule PassthroughModule_16 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_16_io_in),
    .io_out(PassthroughModule_16_io_out)
  );
  PassthroughModule PassthroughModule_17 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_17_io_in),
    .io_out(PassthroughModule_17_io_out)
  );
  PassthroughModule PassthroughModule_18 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_18_io_in),
    .io_out(PassthroughModule_18_io_out)
  );
  PassthroughModule PassthroughModule_19 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_19_io_in),
    .io_out(PassthroughModule_19_io_out)
  );
  PassthroughModule PassthroughModule_20 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_20_io_in),
    .io_out(PassthroughModule_20_io_out)
  );
  PassthroughModule PassthroughModule_21 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_21_io_in),
    .io_out(PassthroughModule_21_io_out)
  );
  PassthroughModule PassthroughModule_22 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_22_io_in),
    .io_out(PassthroughModule_22_io_out)
  );
  PassthroughModule PassthroughModule_23 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_23_io_in),
    .io_out(PassthroughModule_23_io_out)
  );
  PassthroughModule PassthroughModule_24 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_24_io_in),
    .io_out(PassthroughModule_24_io_out)
  );
  PassthroughModule PassthroughModule_25 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_25_io_in),
    .io_out(PassthroughModule_25_io_out)
  );
  PassthroughModule PassthroughModule_26 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_26_io_in),
    .io_out(PassthroughModule_26_io_out)
  );
  PassthroughModule PassthroughModule_27 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_27_io_in),
    .io_out(PassthroughModule_27_io_out)
  );
  PassthroughModule PassthroughModule_28 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_28_io_in),
    .io_out(PassthroughModule_28_io_out)
  );
  PassthroughModule PassthroughModule_29 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_29_io_in),
    .io_out(PassthroughModule_29_io_out)
  );
  PassthroughModule PassthroughModule_30 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_30_io_in),
    .io_out(PassthroughModule_30_io_out)
  );
  PassthroughModule PassthroughModule_31 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_31_io_in),
    .io_out(PassthroughModule_31_io_out)
  );
  PassthroughModule PassthroughModule_32 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_32_io_in),
    .io_out(PassthroughModule_32_io_out)
  );
  PassthroughModule PassthroughModule_33 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_33_io_in),
    .io_out(PassthroughModule_33_io_out)
  );
  PassthroughModule PassthroughModule_34 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_34_io_in),
    .io_out(PassthroughModule_34_io_out)
  );
  PassthroughModule PassthroughModule_35 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_35_io_in),
    .io_out(PassthroughModule_35_io_out)
  );
  PassthroughModule PassthroughModule_36 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_36_io_in),
    .io_out(PassthroughModule_36_io_out)
  );
  PassthroughModule PassthroughModule_37 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_37_io_in),
    .io_out(PassthroughModule_37_io_out)
  );
  PassthroughModule PassthroughModule_38 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_38_io_in),
    .io_out(PassthroughModule_38_io_out)
  );
  PassthroughModule PassthroughModule_39 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_39_io_in),
    .io_out(PassthroughModule_39_io_out)
  );
  PassthroughModule PassthroughModule_40 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_40_io_in),
    .io_out(PassthroughModule_40_io_out)
  );
  PassthroughModule PassthroughModule_41 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_41_io_in),
    .io_out(PassthroughModule_41_io_out)
  );
  PassthroughModule PassthroughModule_42 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_42_io_in),
    .io_out(PassthroughModule_42_io_out)
  );
  PassthroughModule PassthroughModule_43 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_43_io_in),
    .io_out(PassthroughModule_43_io_out)
  );
  PassthroughModule PassthroughModule_44 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_44_io_in),
    .io_out(PassthroughModule_44_io_out)
  );
  PassthroughModule PassthroughModule_45 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_45_io_in),
    .io_out(PassthroughModule_45_io_out)
  );
  PassthroughModule PassthroughModule_46 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_46_io_in),
    .io_out(PassthroughModule_46_io_out)
  );
  PassthroughModule PassthroughModule_47 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_47_io_in),
    .io_out(PassthroughModule_47_io_out)
  );
  PassthroughModule PassthroughModule_48 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_48_io_in),
    .io_out(PassthroughModule_48_io_out)
  );
  PassthroughModule PassthroughModule_49 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_49_io_in),
    .io_out(PassthroughModule_49_io_out)
  );
  PassthroughModule PassthroughModule_50 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_50_io_in),
    .io_out(PassthroughModule_50_io_out)
  );
  PassthroughModule PassthroughModule_51 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_51_io_in),
    .io_out(PassthroughModule_51_io_out)
  );
  PassthroughModule PassthroughModule_52 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_52_io_in),
    .io_out(PassthroughModule_52_io_out)
  );
  PassthroughModule PassthroughModule_53 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_53_io_in),
    .io_out(PassthroughModule_53_io_out)
  );
  PassthroughModule PassthroughModule_54 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_54_io_in),
    .io_out(PassthroughModule_54_io_out)
  );
  PassthroughModule PassthroughModule_55 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_55_io_in),
    .io_out(PassthroughModule_55_io_out)
  );
  PassthroughModule PassthroughModule_56 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_56_io_in),
    .io_out(PassthroughModule_56_io_out)
  );
  PassthroughModule PassthroughModule_57 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_57_io_in),
    .io_out(PassthroughModule_57_io_out)
  );
  PassthroughModule PassthroughModule_58 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_58_io_in),
    .io_out(PassthroughModule_58_io_out)
  );
  PassthroughModule PassthroughModule_59 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_59_io_in),
    .io_out(PassthroughModule_59_io_out)
  );
  PassthroughModule PassthroughModule_60 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_60_io_in),
    .io_out(PassthroughModule_60_io_out)
  );
  PassthroughModule PassthroughModule_61 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_61_io_in),
    .io_out(PassthroughModule_61_io_out)
  );
  PassthroughModule PassthroughModule_62 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_62_io_in),
    .io_out(PassthroughModule_62_io_out)
  );
  PassthroughModule PassthroughModule_63 ( // @[Vec.scala 225:30]
    .io_in(PassthroughModule_63_io_in),
    .io_out(PassthroughModule_63_io_out)
  );
  assign PassthroughModule_io_in = 32'h1; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_1_io_in = 32'h2; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_2_io_in = 32'h3; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_3_io_in = 32'h4; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_4_io_in = 32'h2; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_5_io_in = 32'h3; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_6_io_in = 32'h4; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_7_io_in = 32'h5; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_8_io_in = 32'h3; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_9_io_in = 32'h4; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_10_io_in = 32'h5; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_11_io_in = 32'h6; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_12_io_in = 32'h4; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_13_io_in = 32'h5; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_14_io_in = 32'h6; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_15_io_in = 32'h7; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_16_io_in = 32'h2; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_17_io_in = 32'h3; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_18_io_in = 32'h4; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_19_io_in = 32'h5; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_20_io_in = 32'h3; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_21_io_in = 32'h4; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_22_io_in = 32'h5; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_23_io_in = 32'h6; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_24_io_in = 32'h4; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_25_io_in = 32'h5; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_26_io_in = 32'h6; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_27_io_in = 32'h7; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_28_io_in = 32'h5; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_29_io_in = 32'h6; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_30_io_in = 32'h7; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_31_io_in = 32'h8; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_32_io_in = 32'h3; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_33_io_in = 32'h4; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_34_io_in = 32'h5; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_35_io_in = 32'h6; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_36_io_in = 32'h4; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_37_io_in = 32'h5; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_38_io_in = 32'h6; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_39_io_in = 32'h7; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_40_io_in = 32'h5; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_41_io_in = 32'h6; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_42_io_in = 32'h7; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_43_io_in = 32'h8; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_44_io_in = 32'h6; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_45_io_in = 32'h7; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_46_io_in = 32'h8; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_47_io_in = 32'h9; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_48_io_in = 32'h4; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_49_io_in = 32'h5; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_50_io_in = 32'h6; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_51_io_in = 32'h7; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_52_io_in = 32'h5; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_53_io_in = 32'h6; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_54_io_in = 32'h7; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_55_io_in = 32'h8; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_56_io_in = 32'h6; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_57_io_in = 32'h7; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_58_io_in = 32'h8; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_59_io_in = 32'h9; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_60_io_in = 32'h7; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_61_io_in = 32'h8; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_62_io_in = 32'h9; // @[Vec.scala 217:{43,43}]
  assign PassthroughModule_63_io_in = 32'ha; // @[Vec.scala 217:{43,43}]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_io_out == 32'h1)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_io_out == 32'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_1_io_out == 32'h2)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_1_io_out == 32'h2)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_2_io_out == 32'h3)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_2_io_out == 32'h3)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_3_io_out == 32'h4)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_3_io_out == 32'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_4_io_out == 32'h2)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_4_io_out == 32'h2)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_5_io_out == 32'h3)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_5_io_out == 32'h3)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_6_io_out == 32'h4)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_6_io_out == 32'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_7_io_out == 32'h5)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_7_io_out == 32'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_8_io_out == 32'h3)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_8_io_out == 32'h3)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_9_io_out == 32'h4)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_9_io_out == 32'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_10_io_out == 32'h5)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_10_io_out == 32'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_11_io_out == 32'h6)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_11_io_out == 32'h6)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_12_io_out == 32'h4)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_12_io_out == 32'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_13_io_out == 32'h5)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_13_io_out == 32'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_14_io_out == 32'h6)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_14_io_out == 32'h6)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_15_io_out == 32'h7)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_15_io_out == 32'h7)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_16_io_out == 32'h2)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_16_io_out == 32'h2)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_17_io_out == 32'h3)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_17_io_out == 32'h3)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_18_io_out == 32'h4)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_18_io_out == 32'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_19_io_out == 32'h5)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_19_io_out == 32'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_20_io_out == 32'h3)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_20_io_out == 32'h3)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_21_io_out == 32'h4)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_21_io_out == 32'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_22_io_out == 32'h5)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_22_io_out == 32'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_23_io_out == 32'h6)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_23_io_out == 32'h6)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_24_io_out == 32'h4)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_24_io_out == 32'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_25_io_out == 32'h5)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_25_io_out == 32'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_26_io_out == 32'h6)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_26_io_out == 32'h6)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_27_io_out == 32'h7)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_27_io_out == 32'h7)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_28_io_out == 32'h5)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_28_io_out == 32'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_29_io_out == 32'h6)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_29_io_out == 32'h6)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_30_io_out == 32'h7)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_30_io_out == 32'h7)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_31_io_out == 32'h8)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_31_io_out == 32'h8)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_32_io_out == 32'h3)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_32_io_out == 32'h3)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_33_io_out == 32'h4)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_33_io_out == 32'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_34_io_out == 32'h5)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_34_io_out == 32'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_35_io_out == 32'h6)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_35_io_out == 32'h6)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_36_io_out == 32'h4)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_36_io_out == 32'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_37_io_out == 32'h5)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_37_io_out == 32'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_38_io_out == 32'h6)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_38_io_out == 32'h6)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_39_io_out == 32'h7)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_39_io_out == 32'h7)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_40_io_out == 32'h5)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_40_io_out == 32'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_41_io_out == 32'h6)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_41_io_out == 32'h6)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_42_io_out == 32'h7)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_42_io_out == 32'h7)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_43_io_out == 32'h8)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_43_io_out == 32'h8)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_44_io_out == 32'h6)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_44_io_out == 32'h6)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_45_io_out == 32'h7)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_45_io_out == 32'h7)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_46_io_out == 32'h8)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_46_io_out == 32'h8)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_47_io_out == 32'h9)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_47_io_out == 32'h9)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_48_io_out == 32'h4)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_48_io_out == 32'h4)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_49_io_out == 32'h5)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_49_io_out == 32'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_50_io_out == 32'h6)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_50_io_out == 32'h6)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_51_io_out == 32'h7)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_51_io_out == 32'h7)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_52_io_out == 32'h5)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_52_io_out == 32'h5)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_53_io_out == 32'h6)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_53_io_out == 32'h6)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_54_io_out == 32'h7)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_54_io_out == 32'h7)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_55_io_out == 32'h8)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_55_io_out == 32'h8)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_56_io_out == 32'h6)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_56_io_out == 32'h6)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_57_io_out == 32'h7)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_57_io_out == 32'h7)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_58_io_out == 32'h8)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_58_io_out == 32'h8)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_59_io_out == 32'h9)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_59_io_out == 32'h9)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_60_io_out == 32'h7)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_60_io_out == 32'h7)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_61_io_out == 32'h8)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_61_io_out == 32'h8)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_62_io_out == 32'h9)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_62_io_out == 32'h9)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_63_io_out == 32'ha)) begin
          $fatal; // @[Vec.scala 227:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(PassthroughModule_63_io_out == 32'ha)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Vec.scala:227 assert(receiveMod.out === value.U)\n"); // @[Vec.scala 227:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2) begin
          $finish; // @[Vec.scala 229:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
