module Top(
  input  [7:0] port_foo_bar
);
endmodule
