module IntervalSpec_Anon(
  input   clock,
  input   reset
);
  wire  _T_2 = ~reset; // @[IntervalSpec.scala 878:25]
  wire [6:0] _GEN_0 = 6'sh19 - 6'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_25 = _GEN_0[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [6:0] _GEN_2 = 6'sh1a - 6'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_26 = _GEN_2[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [6:0] _GEN_4 = 6'sh1b - 6'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_27 = _GEN_4[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [6:0] _GEN_6 = 6'sh1c - 6'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_28 = _GEN_6[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [6:0] _GEN_8 = 6'sh1d - 6'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_29 = _GEN_8[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [6:0] _GEN_10 = 6'sh1e - 6'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_30 = _GEN_10[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [6:0] _GEN_12 = 6'sh1f - 6'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_31 = _GEN_12[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [7:0] _GEN_14 = 7'sh20 - 7'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_32 = _GEN_14[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [7:0] _GEN_16 = 7'sh21 - 7'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_33 = _GEN_16[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [7:0] _GEN_18 = 7'sh22 - 7'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_34 = _GEN_18[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [7:0] _GEN_20 = 7'sh23 - 7'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_35 = _GEN_20[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [7:0] _GEN_22 = 7'sh24 - 7'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_36 = _GEN_22[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [7:0] _GEN_24 = 7'sh25 - 7'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_37 = _GEN_24[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [7:0] _GEN_26 = 7'sh26 - 7'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_38 = _GEN_26[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [7:0] _GEN_28 = 7'sh27 - 7'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_39 = _GEN_28[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  wire [7:0] _GEN_30 = 7'sh28 - 7'sh11; // @[IntervalSpec.scala 883:{18,18}]
  wire [5:0] wrappedValue_40 = _GEN_30[5:0]; // @[IntervalSpec.scala 883:{18,18}]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'sh8 == $signed(wrappedValue_25))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'sh8 == $signed(wrappedValue_25))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'sh9 == $signed(wrappedValue_26))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'sh9 == $signed(wrappedValue_26))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'sha == $signed(wrappedValue_27))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'sha == $signed(wrappedValue_27))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'shb == $signed(wrappedValue_28))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'shb == $signed(wrappedValue_28))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'shc == $signed(wrappedValue_29))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'shc == $signed(wrappedValue_29))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'shd == $signed(wrappedValue_30))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'shd == $signed(wrappedValue_30))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'she == $signed(wrappedValue_31))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'she == $signed(wrappedValue_31))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'shf == $signed(wrappedValue_32))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'shf == $signed(wrappedValue_32))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'sh10 == $signed(wrappedValue_33))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'sh10 == $signed(wrappedValue_33))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'sh11 == $signed(wrappedValue_34))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'sh11 == $signed(wrappedValue_34))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'sh12 == $signed(wrappedValue_35))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'sh12 == $signed(wrappedValue_35))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'sh13 == $signed(wrappedValue_36))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'sh13 == $signed(wrappedValue_36))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'sh14 == $signed(wrappedValue_37))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'sh14 == $signed(wrappedValue_37))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'sh15 == $signed(wrappedValue_38))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'sh15 == $signed(wrappedValue_38))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'sh16 == $signed(wrappedValue_39))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'sh16 == $signed(wrappedValue_39))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(6'sh17 == $signed(wrappedValue_40))) begin
          $fatal; // @[IntervalSpec.scala 892:25]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(6'sh17 == $signed(wrappedValue_40))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at IntervalSpec.scala:892 chisel3.assert(goldWrappedValue === wrappedValue)\n"); // @[IntervalSpec.scala 892:25]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2) begin
          $finish; // @[IntervalSpec.scala 895:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
