module M(
  input   clock,
  input   reset
);
  wire  a = 1'h0;
  wire  b_0 = 1'h0;
  wire  b_1 = 1'h0;
endmodule
