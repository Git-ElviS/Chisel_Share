module CastFromNonLit(
  input  [6:0] io_in,
  output [6:0] io_out,
  output       io_valid
);
  assign io_out = io_in; // @[StrongEnum.scala 73:{24,24}]
  assign io_valid = io_out == 7'h0 | io_out == 7'h1 | io_out == 7'h2 | io_out == 7'h64 | io_out == 7'h65; // @[StrongEnum.scala 74:22]
endmodule
module CastFromNonLitTester(
  input   clock,
  input   reset
);
  wire [6:0] mod_io_in; // @[StrongEnum.scala 186:21]
  wire [6:0] mod_io_out; // @[StrongEnum.scala 186:21]
  wire  mod_io_valid; // @[StrongEnum.scala 186:21]
  wire [6:0] mod_1_io_in; // @[StrongEnum.scala 186:21]
  wire [6:0] mod_1_io_out; // @[StrongEnum.scala 186:21]
  wire  mod_1_io_valid; // @[StrongEnum.scala 186:21]
  wire [6:0] mod_2_io_in; // @[StrongEnum.scala 186:21]
  wire [6:0] mod_2_io_out; // @[StrongEnum.scala 186:21]
  wire  mod_2_io_valid; // @[StrongEnum.scala 186:21]
  wire [6:0] mod_3_io_in; // @[StrongEnum.scala 186:21]
  wire [6:0] mod_3_io_out; // @[StrongEnum.scala 186:21]
  wire  mod_3_io_valid; // @[StrongEnum.scala 186:21]
  wire [6:0] mod_4_io_in; // @[StrongEnum.scala 186:21]
  wire [6:0] mod_4_io_out; // @[StrongEnum.scala 186:21]
  wire  mod_4_io_valid; // @[StrongEnum.scala 186:21]
  wire [6:0] mod_5_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_5_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_5_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_6_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_6_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_6_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_7_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_7_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_7_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_8_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_8_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_8_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_9_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_9_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_9_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_10_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_10_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_10_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_11_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_11_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_11_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_12_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_12_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_12_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_13_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_13_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_13_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_14_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_14_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_14_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_15_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_15_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_15_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_16_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_16_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_16_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_17_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_17_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_17_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_18_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_18_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_18_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_19_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_19_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_19_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_20_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_20_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_20_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_21_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_21_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_21_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_22_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_22_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_22_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_23_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_23_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_23_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_24_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_24_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_24_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_25_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_25_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_25_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_26_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_26_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_26_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_27_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_27_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_27_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_28_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_28_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_28_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_29_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_29_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_29_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_30_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_30_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_30_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_31_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_31_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_31_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_32_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_32_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_32_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_33_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_33_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_33_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_34_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_34_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_34_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_35_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_35_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_35_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_36_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_36_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_36_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_37_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_37_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_37_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_38_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_38_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_38_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_39_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_39_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_39_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_40_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_40_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_40_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_41_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_41_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_41_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_42_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_42_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_42_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_43_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_43_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_43_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_44_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_44_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_44_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_45_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_45_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_45_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_46_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_46_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_46_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_47_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_47_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_47_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_48_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_48_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_48_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_49_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_49_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_49_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_50_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_50_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_50_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_51_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_51_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_51_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_52_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_52_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_52_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_53_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_53_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_53_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_54_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_54_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_54_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_55_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_55_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_55_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_56_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_56_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_56_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_57_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_57_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_57_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_58_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_58_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_58_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_59_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_59_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_59_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_60_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_60_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_60_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_61_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_61_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_61_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_62_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_62_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_62_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_63_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_63_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_63_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_64_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_64_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_64_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_65_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_65_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_65_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_66_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_66_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_66_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_67_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_67_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_67_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_68_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_68_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_68_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_69_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_69_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_69_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_70_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_70_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_70_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_71_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_71_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_71_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_72_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_72_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_72_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_73_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_73_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_73_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_74_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_74_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_74_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_75_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_75_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_75_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_76_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_76_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_76_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_77_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_77_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_77_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_78_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_78_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_78_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_79_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_79_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_79_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_80_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_80_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_80_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_81_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_81_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_81_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_82_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_82_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_82_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_83_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_83_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_83_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_84_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_84_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_84_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_85_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_85_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_85_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_86_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_86_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_86_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_87_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_87_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_87_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_88_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_88_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_88_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_89_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_89_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_89_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_90_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_90_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_90_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_91_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_91_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_91_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_92_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_92_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_92_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_93_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_93_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_93_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_94_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_94_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_94_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_95_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_95_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_95_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_96_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_96_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_96_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_97_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_97_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_97_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_98_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_98_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_98_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_99_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_99_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_99_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_100_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_100_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_100_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_101_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_101_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_101_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_102_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_102_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_102_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_103_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_103_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_103_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_104_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_104_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_104_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_105_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_105_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_105_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_106_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_106_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_106_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_107_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_107_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_107_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_108_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_108_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_108_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_109_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_109_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_109_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_110_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_110_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_110_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_111_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_111_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_111_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_112_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_112_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_112_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_113_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_113_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_113_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_114_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_114_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_114_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_115_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_115_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_115_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_116_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_116_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_116_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_117_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_117_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_117_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_118_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_118_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_118_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_119_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_119_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_119_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_120_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_120_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_120_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_121_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_121_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_121_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_122_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_122_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_122_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_123_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_123_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_123_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_124_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_124_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_124_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_125_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_125_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_125_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_126_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_126_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_126_io_valid; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_127_io_in; // @[StrongEnum.scala 196:21]
  wire [6:0] mod_127_io_out; // @[StrongEnum.scala 196:21]
  wire  mod_127_io_valid; // @[StrongEnum.scala 196:21]
  wire  _T_2 = ~reset; // @[StrongEnum.scala 188:11]
  CastFromNonLit mod ( // @[StrongEnum.scala 186:21]
    .io_in(mod_io_in),
    .io_out(mod_io_out),
    .io_valid(mod_io_valid)
  );
  CastFromNonLit mod_1 ( // @[StrongEnum.scala 186:21]
    .io_in(mod_1_io_in),
    .io_out(mod_1_io_out),
    .io_valid(mod_1_io_valid)
  );
  CastFromNonLit mod_2 ( // @[StrongEnum.scala 186:21]
    .io_in(mod_2_io_in),
    .io_out(mod_2_io_out),
    .io_valid(mod_2_io_valid)
  );
  CastFromNonLit mod_3 ( // @[StrongEnum.scala 186:21]
    .io_in(mod_3_io_in),
    .io_out(mod_3_io_out),
    .io_valid(mod_3_io_valid)
  );
  CastFromNonLit mod_4 ( // @[StrongEnum.scala 186:21]
    .io_in(mod_4_io_in),
    .io_out(mod_4_io_out),
    .io_valid(mod_4_io_valid)
  );
  CastFromNonLit mod_5 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_5_io_in),
    .io_out(mod_5_io_out),
    .io_valid(mod_5_io_valid)
  );
  CastFromNonLit mod_6 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_6_io_in),
    .io_out(mod_6_io_out),
    .io_valid(mod_6_io_valid)
  );
  CastFromNonLit mod_7 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_7_io_in),
    .io_out(mod_7_io_out),
    .io_valid(mod_7_io_valid)
  );
  CastFromNonLit mod_8 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_8_io_in),
    .io_out(mod_8_io_out),
    .io_valid(mod_8_io_valid)
  );
  CastFromNonLit mod_9 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_9_io_in),
    .io_out(mod_9_io_out),
    .io_valid(mod_9_io_valid)
  );
  CastFromNonLit mod_10 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_10_io_in),
    .io_out(mod_10_io_out),
    .io_valid(mod_10_io_valid)
  );
  CastFromNonLit mod_11 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_11_io_in),
    .io_out(mod_11_io_out),
    .io_valid(mod_11_io_valid)
  );
  CastFromNonLit mod_12 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_12_io_in),
    .io_out(mod_12_io_out),
    .io_valid(mod_12_io_valid)
  );
  CastFromNonLit mod_13 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_13_io_in),
    .io_out(mod_13_io_out),
    .io_valid(mod_13_io_valid)
  );
  CastFromNonLit mod_14 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_14_io_in),
    .io_out(mod_14_io_out),
    .io_valid(mod_14_io_valid)
  );
  CastFromNonLit mod_15 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_15_io_in),
    .io_out(mod_15_io_out),
    .io_valid(mod_15_io_valid)
  );
  CastFromNonLit mod_16 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_16_io_in),
    .io_out(mod_16_io_out),
    .io_valid(mod_16_io_valid)
  );
  CastFromNonLit mod_17 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_17_io_in),
    .io_out(mod_17_io_out),
    .io_valid(mod_17_io_valid)
  );
  CastFromNonLit mod_18 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_18_io_in),
    .io_out(mod_18_io_out),
    .io_valid(mod_18_io_valid)
  );
  CastFromNonLit mod_19 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_19_io_in),
    .io_out(mod_19_io_out),
    .io_valid(mod_19_io_valid)
  );
  CastFromNonLit mod_20 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_20_io_in),
    .io_out(mod_20_io_out),
    .io_valid(mod_20_io_valid)
  );
  CastFromNonLit mod_21 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_21_io_in),
    .io_out(mod_21_io_out),
    .io_valid(mod_21_io_valid)
  );
  CastFromNonLit mod_22 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_22_io_in),
    .io_out(mod_22_io_out),
    .io_valid(mod_22_io_valid)
  );
  CastFromNonLit mod_23 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_23_io_in),
    .io_out(mod_23_io_out),
    .io_valid(mod_23_io_valid)
  );
  CastFromNonLit mod_24 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_24_io_in),
    .io_out(mod_24_io_out),
    .io_valid(mod_24_io_valid)
  );
  CastFromNonLit mod_25 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_25_io_in),
    .io_out(mod_25_io_out),
    .io_valid(mod_25_io_valid)
  );
  CastFromNonLit mod_26 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_26_io_in),
    .io_out(mod_26_io_out),
    .io_valid(mod_26_io_valid)
  );
  CastFromNonLit mod_27 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_27_io_in),
    .io_out(mod_27_io_out),
    .io_valid(mod_27_io_valid)
  );
  CastFromNonLit mod_28 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_28_io_in),
    .io_out(mod_28_io_out),
    .io_valid(mod_28_io_valid)
  );
  CastFromNonLit mod_29 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_29_io_in),
    .io_out(mod_29_io_out),
    .io_valid(mod_29_io_valid)
  );
  CastFromNonLit mod_30 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_30_io_in),
    .io_out(mod_30_io_out),
    .io_valid(mod_30_io_valid)
  );
  CastFromNonLit mod_31 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_31_io_in),
    .io_out(mod_31_io_out),
    .io_valid(mod_31_io_valid)
  );
  CastFromNonLit mod_32 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_32_io_in),
    .io_out(mod_32_io_out),
    .io_valid(mod_32_io_valid)
  );
  CastFromNonLit mod_33 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_33_io_in),
    .io_out(mod_33_io_out),
    .io_valid(mod_33_io_valid)
  );
  CastFromNonLit mod_34 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_34_io_in),
    .io_out(mod_34_io_out),
    .io_valid(mod_34_io_valid)
  );
  CastFromNonLit mod_35 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_35_io_in),
    .io_out(mod_35_io_out),
    .io_valid(mod_35_io_valid)
  );
  CastFromNonLit mod_36 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_36_io_in),
    .io_out(mod_36_io_out),
    .io_valid(mod_36_io_valid)
  );
  CastFromNonLit mod_37 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_37_io_in),
    .io_out(mod_37_io_out),
    .io_valid(mod_37_io_valid)
  );
  CastFromNonLit mod_38 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_38_io_in),
    .io_out(mod_38_io_out),
    .io_valid(mod_38_io_valid)
  );
  CastFromNonLit mod_39 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_39_io_in),
    .io_out(mod_39_io_out),
    .io_valid(mod_39_io_valid)
  );
  CastFromNonLit mod_40 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_40_io_in),
    .io_out(mod_40_io_out),
    .io_valid(mod_40_io_valid)
  );
  CastFromNonLit mod_41 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_41_io_in),
    .io_out(mod_41_io_out),
    .io_valid(mod_41_io_valid)
  );
  CastFromNonLit mod_42 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_42_io_in),
    .io_out(mod_42_io_out),
    .io_valid(mod_42_io_valid)
  );
  CastFromNonLit mod_43 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_43_io_in),
    .io_out(mod_43_io_out),
    .io_valid(mod_43_io_valid)
  );
  CastFromNonLit mod_44 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_44_io_in),
    .io_out(mod_44_io_out),
    .io_valid(mod_44_io_valid)
  );
  CastFromNonLit mod_45 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_45_io_in),
    .io_out(mod_45_io_out),
    .io_valid(mod_45_io_valid)
  );
  CastFromNonLit mod_46 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_46_io_in),
    .io_out(mod_46_io_out),
    .io_valid(mod_46_io_valid)
  );
  CastFromNonLit mod_47 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_47_io_in),
    .io_out(mod_47_io_out),
    .io_valid(mod_47_io_valid)
  );
  CastFromNonLit mod_48 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_48_io_in),
    .io_out(mod_48_io_out),
    .io_valid(mod_48_io_valid)
  );
  CastFromNonLit mod_49 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_49_io_in),
    .io_out(mod_49_io_out),
    .io_valid(mod_49_io_valid)
  );
  CastFromNonLit mod_50 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_50_io_in),
    .io_out(mod_50_io_out),
    .io_valid(mod_50_io_valid)
  );
  CastFromNonLit mod_51 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_51_io_in),
    .io_out(mod_51_io_out),
    .io_valid(mod_51_io_valid)
  );
  CastFromNonLit mod_52 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_52_io_in),
    .io_out(mod_52_io_out),
    .io_valid(mod_52_io_valid)
  );
  CastFromNonLit mod_53 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_53_io_in),
    .io_out(mod_53_io_out),
    .io_valid(mod_53_io_valid)
  );
  CastFromNonLit mod_54 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_54_io_in),
    .io_out(mod_54_io_out),
    .io_valid(mod_54_io_valid)
  );
  CastFromNonLit mod_55 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_55_io_in),
    .io_out(mod_55_io_out),
    .io_valid(mod_55_io_valid)
  );
  CastFromNonLit mod_56 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_56_io_in),
    .io_out(mod_56_io_out),
    .io_valid(mod_56_io_valid)
  );
  CastFromNonLit mod_57 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_57_io_in),
    .io_out(mod_57_io_out),
    .io_valid(mod_57_io_valid)
  );
  CastFromNonLit mod_58 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_58_io_in),
    .io_out(mod_58_io_out),
    .io_valid(mod_58_io_valid)
  );
  CastFromNonLit mod_59 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_59_io_in),
    .io_out(mod_59_io_out),
    .io_valid(mod_59_io_valid)
  );
  CastFromNonLit mod_60 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_60_io_in),
    .io_out(mod_60_io_out),
    .io_valid(mod_60_io_valid)
  );
  CastFromNonLit mod_61 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_61_io_in),
    .io_out(mod_61_io_out),
    .io_valid(mod_61_io_valid)
  );
  CastFromNonLit mod_62 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_62_io_in),
    .io_out(mod_62_io_out),
    .io_valid(mod_62_io_valid)
  );
  CastFromNonLit mod_63 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_63_io_in),
    .io_out(mod_63_io_out),
    .io_valid(mod_63_io_valid)
  );
  CastFromNonLit mod_64 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_64_io_in),
    .io_out(mod_64_io_out),
    .io_valid(mod_64_io_valid)
  );
  CastFromNonLit mod_65 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_65_io_in),
    .io_out(mod_65_io_out),
    .io_valid(mod_65_io_valid)
  );
  CastFromNonLit mod_66 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_66_io_in),
    .io_out(mod_66_io_out),
    .io_valid(mod_66_io_valid)
  );
  CastFromNonLit mod_67 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_67_io_in),
    .io_out(mod_67_io_out),
    .io_valid(mod_67_io_valid)
  );
  CastFromNonLit mod_68 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_68_io_in),
    .io_out(mod_68_io_out),
    .io_valid(mod_68_io_valid)
  );
  CastFromNonLit mod_69 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_69_io_in),
    .io_out(mod_69_io_out),
    .io_valid(mod_69_io_valid)
  );
  CastFromNonLit mod_70 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_70_io_in),
    .io_out(mod_70_io_out),
    .io_valid(mod_70_io_valid)
  );
  CastFromNonLit mod_71 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_71_io_in),
    .io_out(mod_71_io_out),
    .io_valid(mod_71_io_valid)
  );
  CastFromNonLit mod_72 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_72_io_in),
    .io_out(mod_72_io_out),
    .io_valid(mod_72_io_valid)
  );
  CastFromNonLit mod_73 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_73_io_in),
    .io_out(mod_73_io_out),
    .io_valid(mod_73_io_valid)
  );
  CastFromNonLit mod_74 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_74_io_in),
    .io_out(mod_74_io_out),
    .io_valid(mod_74_io_valid)
  );
  CastFromNonLit mod_75 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_75_io_in),
    .io_out(mod_75_io_out),
    .io_valid(mod_75_io_valid)
  );
  CastFromNonLit mod_76 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_76_io_in),
    .io_out(mod_76_io_out),
    .io_valid(mod_76_io_valid)
  );
  CastFromNonLit mod_77 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_77_io_in),
    .io_out(mod_77_io_out),
    .io_valid(mod_77_io_valid)
  );
  CastFromNonLit mod_78 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_78_io_in),
    .io_out(mod_78_io_out),
    .io_valid(mod_78_io_valid)
  );
  CastFromNonLit mod_79 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_79_io_in),
    .io_out(mod_79_io_out),
    .io_valid(mod_79_io_valid)
  );
  CastFromNonLit mod_80 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_80_io_in),
    .io_out(mod_80_io_out),
    .io_valid(mod_80_io_valid)
  );
  CastFromNonLit mod_81 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_81_io_in),
    .io_out(mod_81_io_out),
    .io_valid(mod_81_io_valid)
  );
  CastFromNonLit mod_82 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_82_io_in),
    .io_out(mod_82_io_out),
    .io_valid(mod_82_io_valid)
  );
  CastFromNonLit mod_83 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_83_io_in),
    .io_out(mod_83_io_out),
    .io_valid(mod_83_io_valid)
  );
  CastFromNonLit mod_84 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_84_io_in),
    .io_out(mod_84_io_out),
    .io_valid(mod_84_io_valid)
  );
  CastFromNonLit mod_85 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_85_io_in),
    .io_out(mod_85_io_out),
    .io_valid(mod_85_io_valid)
  );
  CastFromNonLit mod_86 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_86_io_in),
    .io_out(mod_86_io_out),
    .io_valid(mod_86_io_valid)
  );
  CastFromNonLit mod_87 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_87_io_in),
    .io_out(mod_87_io_out),
    .io_valid(mod_87_io_valid)
  );
  CastFromNonLit mod_88 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_88_io_in),
    .io_out(mod_88_io_out),
    .io_valid(mod_88_io_valid)
  );
  CastFromNonLit mod_89 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_89_io_in),
    .io_out(mod_89_io_out),
    .io_valid(mod_89_io_valid)
  );
  CastFromNonLit mod_90 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_90_io_in),
    .io_out(mod_90_io_out),
    .io_valid(mod_90_io_valid)
  );
  CastFromNonLit mod_91 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_91_io_in),
    .io_out(mod_91_io_out),
    .io_valid(mod_91_io_valid)
  );
  CastFromNonLit mod_92 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_92_io_in),
    .io_out(mod_92_io_out),
    .io_valid(mod_92_io_valid)
  );
  CastFromNonLit mod_93 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_93_io_in),
    .io_out(mod_93_io_out),
    .io_valid(mod_93_io_valid)
  );
  CastFromNonLit mod_94 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_94_io_in),
    .io_out(mod_94_io_out),
    .io_valid(mod_94_io_valid)
  );
  CastFromNonLit mod_95 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_95_io_in),
    .io_out(mod_95_io_out),
    .io_valid(mod_95_io_valid)
  );
  CastFromNonLit mod_96 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_96_io_in),
    .io_out(mod_96_io_out),
    .io_valid(mod_96_io_valid)
  );
  CastFromNonLit mod_97 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_97_io_in),
    .io_out(mod_97_io_out),
    .io_valid(mod_97_io_valid)
  );
  CastFromNonLit mod_98 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_98_io_in),
    .io_out(mod_98_io_out),
    .io_valid(mod_98_io_valid)
  );
  CastFromNonLit mod_99 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_99_io_in),
    .io_out(mod_99_io_out),
    .io_valid(mod_99_io_valid)
  );
  CastFromNonLit mod_100 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_100_io_in),
    .io_out(mod_100_io_out),
    .io_valid(mod_100_io_valid)
  );
  CastFromNonLit mod_101 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_101_io_in),
    .io_out(mod_101_io_out),
    .io_valid(mod_101_io_valid)
  );
  CastFromNonLit mod_102 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_102_io_in),
    .io_out(mod_102_io_out),
    .io_valid(mod_102_io_valid)
  );
  CastFromNonLit mod_103 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_103_io_in),
    .io_out(mod_103_io_out),
    .io_valid(mod_103_io_valid)
  );
  CastFromNonLit mod_104 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_104_io_in),
    .io_out(mod_104_io_out),
    .io_valid(mod_104_io_valid)
  );
  CastFromNonLit mod_105 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_105_io_in),
    .io_out(mod_105_io_out),
    .io_valid(mod_105_io_valid)
  );
  CastFromNonLit mod_106 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_106_io_in),
    .io_out(mod_106_io_out),
    .io_valid(mod_106_io_valid)
  );
  CastFromNonLit mod_107 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_107_io_in),
    .io_out(mod_107_io_out),
    .io_valid(mod_107_io_valid)
  );
  CastFromNonLit mod_108 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_108_io_in),
    .io_out(mod_108_io_out),
    .io_valid(mod_108_io_valid)
  );
  CastFromNonLit mod_109 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_109_io_in),
    .io_out(mod_109_io_out),
    .io_valid(mod_109_io_valid)
  );
  CastFromNonLit mod_110 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_110_io_in),
    .io_out(mod_110_io_out),
    .io_valid(mod_110_io_valid)
  );
  CastFromNonLit mod_111 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_111_io_in),
    .io_out(mod_111_io_out),
    .io_valid(mod_111_io_valid)
  );
  CastFromNonLit mod_112 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_112_io_in),
    .io_out(mod_112_io_out),
    .io_valid(mod_112_io_valid)
  );
  CastFromNonLit mod_113 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_113_io_in),
    .io_out(mod_113_io_out),
    .io_valid(mod_113_io_valid)
  );
  CastFromNonLit mod_114 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_114_io_in),
    .io_out(mod_114_io_out),
    .io_valid(mod_114_io_valid)
  );
  CastFromNonLit mod_115 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_115_io_in),
    .io_out(mod_115_io_out),
    .io_valid(mod_115_io_valid)
  );
  CastFromNonLit mod_116 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_116_io_in),
    .io_out(mod_116_io_out),
    .io_valid(mod_116_io_valid)
  );
  CastFromNonLit mod_117 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_117_io_in),
    .io_out(mod_117_io_out),
    .io_valid(mod_117_io_valid)
  );
  CastFromNonLit mod_118 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_118_io_in),
    .io_out(mod_118_io_out),
    .io_valid(mod_118_io_valid)
  );
  CastFromNonLit mod_119 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_119_io_in),
    .io_out(mod_119_io_out),
    .io_valid(mod_119_io_valid)
  );
  CastFromNonLit mod_120 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_120_io_in),
    .io_out(mod_120_io_out),
    .io_valid(mod_120_io_valid)
  );
  CastFromNonLit mod_121 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_121_io_in),
    .io_out(mod_121_io_out),
    .io_valid(mod_121_io_valid)
  );
  CastFromNonLit mod_122 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_122_io_in),
    .io_out(mod_122_io_out),
    .io_valid(mod_122_io_valid)
  );
  CastFromNonLit mod_123 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_123_io_in),
    .io_out(mod_123_io_out),
    .io_valid(mod_123_io_valid)
  );
  CastFromNonLit mod_124 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_124_io_in),
    .io_out(mod_124_io_out),
    .io_valid(mod_124_io_valid)
  );
  CastFromNonLit mod_125 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_125_io_in),
    .io_out(mod_125_io_out),
    .io_valid(mod_125_io_valid)
  );
  CastFromNonLit mod_126 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_126_io_in),
    .io_out(mod_126_io_out),
    .io_valid(mod_126_io_valid)
  );
  CastFromNonLit mod_127 ( // @[StrongEnum.scala 196:21]
    .io_in(mod_127_io_in),
    .io_out(mod_127_io_out),
    .io_valid(mod_127_io_valid)
  );
  assign mod_io_in = 7'h0; // @[StrongEnum.scala 187:15]
  assign mod_1_io_in = 7'h1; // @[StrongEnum.scala 187:15]
  assign mod_2_io_in = 7'h2; // @[StrongEnum.scala 187:15]
  assign mod_3_io_in = 7'h64; // @[StrongEnum.scala 187:15]
  assign mod_4_io_in = 7'h65; // @[StrongEnum.scala 187:15]
  assign mod_5_io_in = 7'h3; // @[StrongEnum.scala 197:15]
  assign mod_6_io_in = 7'h4; // @[StrongEnum.scala 197:15]
  assign mod_7_io_in = 7'h5; // @[StrongEnum.scala 197:15]
  assign mod_8_io_in = 7'h6; // @[StrongEnum.scala 197:15]
  assign mod_9_io_in = 7'h7; // @[StrongEnum.scala 197:15]
  assign mod_10_io_in = 7'h8; // @[StrongEnum.scala 197:15]
  assign mod_11_io_in = 7'h9; // @[StrongEnum.scala 197:15]
  assign mod_12_io_in = 7'ha; // @[StrongEnum.scala 197:15]
  assign mod_13_io_in = 7'hb; // @[StrongEnum.scala 197:15]
  assign mod_14_io_in = 7'hc; // @[StrongEnum.scala 197:15]
  assign mod_15_io_in = 7'hd; // @[StrongEnum.scala 197:15]
  assign mod_16_io_in = 7'he; // @[StrongEnum.scala 197:15]
  assign mod_17_io_in = 7'hf; // @[StrongEnum.scala 197:15]
  assign mod_18_io_in = 7'h10; // @[StrongEnum.scala 197:15]
  assign mod_19_io_in = 7'h11; // @[StrongEnum.scala 197:15]
  assign mod_20_io_in = 7'h12; // @[StrongEnum.scala 197:15]
  assign mod_21_io_in = 7'h13; // @[StrongEnum.scala 197:15]
  assign mod_22_io_in = 7'h14; // @[StrongEnum.scala 197:15]
  assign mod_23_io_in = 7'h15; // @[StrongEnum.scala 197:15]
  assign mod_24_io_in = 7'h16; // @[StrongEnum.scala 197:15]
  assign mod_25_io_in = 7'h17; // @[StrongEnum.scala 197:15]
  assign mod_26_io_in = 7'h18; // @[StrongEnum.scala 197:15]
  assign mod_27_io_in = 7'h19; // @[StrongEnum.scala 197:15]
  assign mod_28_io_in = 7'h1a; // @[StrongEnum.scala 197:15]
  assign mod_29_io_in = 7'h1b; // @[StrongEnum.scala 197:15]
  assign mod_30_io_in = 7'h1c; // @[StrongEnum.scala 197:15]
  assign mod_31_io_in = 7'h1d; // @[StrongEnum.scala 197:15]
  assign mod_32_io_in = 7'h1e; // @[StrongEnum.scala 197:15]
  assign mod_33_io_in = 7'h1f; // @[StrongEnum.scala 197:15]
  assign mod_34_io_in = 7'h20; // @[StrongEnum.scala 197:15]
  assign mod_35_io_in = 7'h21; // @[StrongEnum.scala 197:15]
  assign mod_36_io_in = 7'h22; // @[StrongEnum.scala 197:15]
  assign mod_37_io_in = 7'h23; // @[StrongEnum.scala 197:15]
  assign mod_38_io_in = 7'h24; // @[StrongEnum.scala 197:15]
  assign mod_39_io_in = 7'h25; // @[StrongEnum.scala 197:15]
  assign mod_40_io_in = 7'h26; // @[StrongEnum.scala 197:15]
  assign mod_41_io_in = 7'h27; // @[StrongEnum.scala 197:15]
  assign mod_42_io_in = 7'h28; // @[StrongEnum.scala 197:15]
  assign mod_43_io_in = 7'h29; // @[StrongEnum.scala 197:15]
  assign mod_44_io_in = 7'h2a; // @[StrongEnum.scala 197:15]
  assign mod_45_io_in = 7'h2b; // @[StrongEnum.scala 197:15]
  assign mod_46_io_in = 7'h2c; // @[StrongEnum.scala 197:15]
  assign mod_47_io_in = 7'h2d; // @[StrongEnum.scala 197:15]
  assign mod_48_io_in = 7'h2e; // @[StrongEnum.scala 197:15]
  assign mod_49_io_in = 7'h2f; // @[StrongEnum.scala 197:15]
  assign mod_50_io_in = 7'h30; // @[StrongEnum.scala 197:15]
  assign mod_51_io_in = 7'h31; // @[StrongEnum.scala 197:15]
  assign mod_52_io_in = 7'h32; // @[StrongEnum.scala 197:15]
  assign mod_53_io_in = 7'h33; // @[StrongEnum.scala 197:15]
  assign mod_54_io_in = 7'h34; // @[StrongEnum.scala 197:15]
  assign mod_55_io_in = 7'h35; // @[StrongEnum.scala 197:15]
  assign mod_56_io_in = 7'h36; // @[StrongEnum.scala 197:15]
  assign mod_57_io_in = 7'h37; // @[StrongEnum.scala 197:15]
  assign mod_58_io_in = 7'h38; // @[StrongEnum.scala 197:15]
  assign mod_59_io_in = 7'h39; // @[StrongEnum.scala 197:15]
  assign mod_60_io_in = 7'h3a; // @[StrongEnum.scala 197:15]
  assign mod_61_io_in = 7'h3b; // @[StrongEnum.scala 197:15]
  assign mod_62_io_in = 7'h3c; // @[StrongEnum.scala 197:15]
  assign mod_63_io_in = 7'h3d; // @[StrongEnum.scala 197:15]
  assign mod_64_io_in = 7'h3e; // @[StrongEnum.scala 197:15]
  assign mod_65_io_in = 7'h3f; // @[StrongEnum.scala 197:15]
  assign mod_66_io_in = 7'h40; // @[StrongEnum.scala 197:15]
  assign mod_67_io_in = 7'h41; // @[StrongEnum.scala 197:15]
  assign mod_68_io_in = 7'h42; // @[StrongEnum.scala 197:15]
  assign mod_69_io_in = 7'h43; // @[StrongEnum.scala 197:15]
  assign mod_70_io_in = 7'h44; // @[StrongEnum.scala 197:15]
  assign mod_71_io_in = 7'h45; // @[StrongEnum.scala 197:15]
  assign mod_72_io_in = 7'h46; // @[StrongEnum.scala 197:15]
  assign mod_73_io_in = 7'h47; // @[StrongEnum.scala 197:15]
  assign mod_74_io_in = 7'h48; // @[StrongEnum.scala 197:15]
  assign mod_75_io_in = 7'h49; // @[StrongEnum.scala 197:15]
  assign mod_76_io_in = 7'h4a; // @[StrongEnum.scala 197:15]
  assign mod_77_io_in = 7'h4b; // @[StrongEnum.scala 197:15]
  assign mod_78_io_in = 7'h4c; // @[StrongEnum.scala 197:15]
  assign mod_79_io_in = 7'h4d; // @[StrongEnum.scala 197:15]
  assign mod_80_io_in = 7'h4e; // @[StrongEnum.scala 197:15]
  assign mod_81_io_in = 7'h4f; // @[StrongEnum.scala 197:15]
  assign mod_82_io_in = 7'h50; // @[StrongEnum.scala 197:15]
  assign mod_83_io_in = 7'h51; // @[StrongEnum.scala 197:15]
  assign mod_84_io_in = 7'h52; // @[StrongEnum.scala 197:15]
  assign mod_85_io_in = 7'h53; // @[StrongEnum.scala 197:15]
  assign mod_86_io_in = 7'h54; // @[StrongEnum.scala 197:15]
  assign mod_87_io_in = 7'h55; // @[StrongEnum.scala 197:15]
  assign mod_88_io_in = 7'h56; // @[StrongEnum.scala 197:15]
  assign mod_89_io_in = 7'h57; // @[StrongEnum.scala 197:15]
  assign mod_90_io_in = 7'h58; // @[StrongEnum.scala 197:15]
  assign mod_91_io_in = 7'h59; // @[StrongEnum.scala 197:15]
  assign mod_92_io_in = 7'h5a; // @[StrongEnum.scala 197:15]
  assign mod_93_io_in = 7'h5b; // @[StrongEnum.scala 197:15]
  assign mod_94_io_in = 7'h5c; // @[StrongEnum.scala 197:15]
  assign mod_95_io_in = 7'h5d; // @[StrongEnum.scala 197:15]
  assign mod_96_io_in = 7'h5e; // @[StrongEnum.scala 197:15]
  assign mod_97_io_in = 7'h5f; // @[StrongEnum.scala 197:15]
  assign mod_98_io_in = 7'h60; // @[StrongEnum.scala 197:15]
  assign mod_99_io_in = 7'h61; // @[StrongEnum.scala 197:15]
  assign mod_100_io_in = 7'h62; // @[StrongEnum.scala 197:15]
  assign mod_101_io_in = 7'h63; // @[StrongEnum.scala 197:15]
  assign mod_102_io_in = 7'h66; // @[StrongEnum.scala 197:15]
  assign mod_103_io_in = 7'h67; // @[StrongEnum.scala 197:15]
  assign mod_104_io_in = 7'h68; // @[StrongEnum.scala 197:15]
  assign mod_105_io_in = 7'h69; // @[StrongEnum.scala 197:15]
  assign mod_106_io_in = 7'h6a; // @[StrongEnum.scala 197:15]
  assign mod_107_io_in = 7'h6b; // @[StrongEnum.scala 197:15]
  assign mod_108_io_in = 7'h6c; // @[StrongEnum.scala 197:15]
  assign mod_109_io_in = 7'h6d; // @[StrongEnum.scala 197:15]
  assign mod_110_io_in = 7'h6e; // @[StrongEnum.scala 197:15]
  assign mod_111_io_in = 7'h6f; // @[StrongEnum.scala 197:15]
  assign mod_112_io_in = 7'h70; // @[StrongEnum.scala 197:15]
  assign mod_113_io_in = 7'h71; // @[StrongEnum.scala 197:15]
  assign mod_114_io_in = 7'h72; // @[StrongEnum.scala 197:15]
  assign mod_115_io_in = 7'h73; // @[StrongEnum.scala 197:15]
  assign mod_116_io_in = 7'h74; // @[StrongEnum.scala 197:15]
  assign mod_117_io_in = 7'h75; // @[StrongEnum.scala 197:15]
  assign mod_118_io_in = 7'h76; // @[StrongEnum.scala 197:15]
  assign mod_119_io_in = 7'h77; // @[StrongEnum.scala 197:15]
  assign mod_120_io_in = 7'h78; // @[StrongEnum.scala 197:15]
  assign mod_121_io_in = 7'h79; // @[StrongEnum.scala 197:15]
  assign mod_122_io_in = 7'h7a; // @[StrongEnum.scala 197:15]
  assign mod_123_io_in = 7'h7b; // @[StrongEnum.scala 197:15]
  assign mod_124_io_in = 7'h7c; // @[StrongEnum.scala 197:15]
  assign mod_125_io_in = 7'h7d; // @[StrongEnum.scala 197:15]
  assign mod_126_io_in = 7'h7e; // @[StrongEnum.scala 197:15]
  assign mod_127_io_in = 7'h7f; // @[StrongEnum.scala 197:15]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(mod_io_out == 7'h0)) begin
          $fatal; // @[StrongEnum.scala 188:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(mod_io_out == 7'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:188 assert(mod.io.out === enum)\n"); // @[StrongEnum.scala 188:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~mod_io_valid) begin
          $fatal; // @[StrongEnum.scala 189:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~mod_io_valid) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:189 assert(mod.io.valid === true.B)\n"); // @[StrongEnum.scala 189:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(mod_1_io_out == 7'h1)) begin
          $fatal; // @[StrongEnum.scala 188:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(mod_1_io_out == 7'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:188 assert(mod.io.out === enum)\n"); // @[StrongEnum.scala 188:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~mod_1_io_valid) begin
          $fatal; // @[StrongEnum.scala 189:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~mod_1_io_valid) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:189 assert(mod.io.valid === true.B)\n"); // @[StrongEnum.scala 189:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(mod_2_io_out == 7'h2)) begin
          $fatal; // @[StrongEnum.scala 188:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(mod_2_io_out == 7'h2)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:188 assert(mod.io.out === enum)\n"); // @[StrongEnum.scala 188:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~mod_2_io_valid) begin
          $fatal; // @[StrongEnum.scala 189:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~mod_2_io_valid) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:189 assert(mod.io.valid === true.B)\n"); // @[StrongEnum.scala 189:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(mod_3_io_out == 7'h64)) begin
          $fatal; // @[StrongEnum.scala 188:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(mod_3_io_out == 7'h64)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:188 assert(mod.io.out === enum)\n"); // @[StrongEnum.scala 188:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~mod_3_io_valid) begin
          $fatal; // @[StrongEnum.scala 189:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~mod_3_io_valid) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:189 assert(mod.io.valid === true.B)\n"); // @[StrongEnum.scala 189:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(mod_4_io_out == 7'h65)) begin
          $fatal; // @[StrongEnum.scala 188:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(mod_4_io_out == 7'h65)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:188 assert(mod.io.out === enum)\n"); // @[StrongEnum.scala 188:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~mod_4_io_valid) begin
          $fatal; // @[StrongEnum.scala 189:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~mod_4_io_valid) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:189 assert(mod.io.valid === true.B)\n"); // @[StrongEnum.scala 189:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_5_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_5_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_6_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_6_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_7_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_7_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_8_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_8_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_9_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_9_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_10_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_10_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_11_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_11_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_12_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_12_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_13_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_13_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_14_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_14_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_15_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_15_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_16_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_16_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_17_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_17_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_18_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_18_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_19_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_19_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_20_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_20_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_21_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_21_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_22_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_22_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_23_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_23_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_24_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_24_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_25_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_25_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_26_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_26_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_27_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_27_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_28_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_28_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_29_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_29_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_30_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_30_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_31_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_31_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_32_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_32_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_33_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_33_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_34_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_34_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_35_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_35_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_36_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_36_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_37_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_37_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_38_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_38_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_39_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_39_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_40_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_40_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_41_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_41_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_42_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_42_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_43_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_43_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_44_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_44_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_45_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_45_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_46_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_46_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_47_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_47_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_48_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_48_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_49_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_49_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_50_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_50_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_51_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_51_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_52_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_52_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_53_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_53_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_54_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_54_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_55_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_55_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_56_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_56_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_57_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_57_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_58_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_58_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_59_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_59_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_60_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_60_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_61_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_61_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_62_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_62_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_63_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_63_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_64_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_64_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_65_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_65_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_66_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_66_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_67_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_67_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_68_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_68_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_69_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_69_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_70_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_70_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_71_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_71_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_72_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_72_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_73_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_73_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_74_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_74_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_75_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_75_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_76_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_76_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_77_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_77_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_78_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_78_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_79_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_79_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_80_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_80_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_81_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_81_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_82_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_82_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_83_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_83_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_84_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_84_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_85_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_85_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_86_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_86_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_87_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_87_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_88_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_88_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_89_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_89_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_90_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_90_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_91_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_91_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_92_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_92_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_93_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_93_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_94_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_94_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_95_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_95_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_96_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_96_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_97_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_97_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_98_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_98_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_99_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_99_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_100_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_100_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_101_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_101_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_102_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_102_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_103_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_103_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_104_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_104_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_105_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_105_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_106_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_106_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_107_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_107_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_108_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_108_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_109_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_109_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_110_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_110_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_111_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_111_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_112_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_112_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_113_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_113_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_114_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_114_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_115_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_115_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_116_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_116_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_117_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_117_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_118_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_118_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_119_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_119_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_120_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_120_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_121_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_121_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_122_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_122_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_123_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_123_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_124_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_124_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_125_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_125_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_126_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_126_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(~mod_127_io_valid)) begin
          $fatal; // @[StrongEnum.scala 199:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(~mod_127_io_valid)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at StrongEnum.scala:199 assert(mod.io.valid === false.B)\n"); // @[StrongEnum.scala 199:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2) begin
          $finish; // @[StrongEnum.scala 202:7]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
